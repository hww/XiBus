module ntc (
	input clk,    // Clock
	input rst_n,  // Asynchronous reset active low
	inout ad[31:0],	// Address Data Bus
);

ic74als651(
	);

endmodule : ntc